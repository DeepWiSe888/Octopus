
module global_clk (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
